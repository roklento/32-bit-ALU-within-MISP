module myOr(
output [31:0] R,
input [31:0] A,
input [31:0] B
);

	or (R[0],A[0],B[0]);
	or (R[1],A[1],B[1]);
	or (R[2],A[2],B[2]);
	or (R[3],A[3],B[3]);
	or (R[4],A[4],B[4]);
	or (R[5],A[5],B[5]);
	or (R[6],A[6],B[6]);
	or (R[7],A[7],B[7]);
	or (R[8],A[8],B[8]);
	or (R[9],A[9],B[9]);
	or (R[10],A[10],B[10]);
	or (R[11],A[11],B[11]);
	or (R[12],A[12],B[12]);
	or (R[13],A[13],B[13]);
	or (R[14],A[14],B[14]);
	or (R[15],A[15],B[15]);
	or (R[16],A[16],B[16]);
	or (R[17],A[17],B[17]);
	or (R[18],A[18],B[18]);
	or (R[19],A[19],B[19]);
	or (R[20],A[20],B[20]);
	or (R[21],A[21],B[21]);
	or (R[22],A[22],B[22]);
	or (R[23],A[23],B[23]);
	or (R[24],A[24],B[24]);
	or (R[25],A[25],B[25]);
	or (R[26],A[26],B[26]);
	or (R[27],A[27],B[27]);
	or (R[28],A[28],B[28]);
	or (R[29],A[29],B[29]);
	or (R[30],A[30],B[30]);
	or (R[31],A[31],B[31]);



endmodule